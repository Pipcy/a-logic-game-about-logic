`timescale 1ns / 1ps

module player_controller_tb(

    );
endmodule
